`timescale 1ns/1ps

module TopTop_tb;

//parameter SIZE = 1;
parameter[15:0] SIZE = 16'h0202;
parameter MAX_WORD_LENGTH = 32;

//inputs
reg clk, reset, start;
reg[31:0] instruction;
//reg[5:0] LENGTH;



reg external;
reg[7:0] Tile_i = 8'b0;
reg[7:0] Tile_j = 8'b0;
reg[7:0] BRAM_i = 8'b0;
reg[7:0] BRAM_j = 8'b0;
reg WEA, WEB, mode;
reg[9:0] ADDRA = -1;
reg[9:0] ADDRB = 5;
reg[15:0] DINA, DINB;
wire[15:0] DOUTA, DOUTB;
reg[159:0] ram[15:0];
reg[9:0] ram_ptr = 0;
reg[1:0] Activation_Function;
reg Tanh_In;
integer i=0, j=0, k=0;
// reg[0:4*SIZE*MAX_WORD_LENGTH-1] EAST_I;
// reg[0:4*SIZE*MAX_WORD_LENGTH-1] WEST_I;
// wire[0:4*SIZE*MAX_WORD_LENGTH-1] Y;

TopTop #(SIZE[15:8], SIZE[7:0], MAX_WORD_LENGTH) TopTopTB(clk, reset, start, instruction, external, Tile_i, Tile_j, BRAM_i, BRAM_j, WEA, 1'b0, ADDRA, ADDRB, DINA, DINB, DOUTA, DOUTB, Activation_Function, Tanh_In);

initial begin
  clk = 1;
  forever #5 clk = !clk;
end

always @ (posedge clk) begin

    // for(i=0; i<1; i=i+1) begin
    //     for(j=0; j<1; j=j+1) begin
           
    //     end
    // end
    if(Tile_i == 0 && Tile_j == 0 && BRAM_i == 0 && BRAM_j == 0) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
           
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
	if(Tile_i == 0 && Tile_j == 0 && BRAM_i == 0 && BRAM_j == 1) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
            
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
    if(Tile_i == 0 && Tile_j == 0 && BRAM_i == 1 && BRAM_j == 0) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
           
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
    if(Tile_i == 0 && Tile_j == 0 && BRAM_i == 1 && BRAM_j == 1) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
           
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
	
	
	if(Tile_i == 0 && Tile_j == 1 && BRAM_i == 0 && BRAM_j == 0) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
           
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
    if(Tile_i == 0 && Tile_j == 1 && BRAM_i == 0 && BRAM_j == 1) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
            
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
    if(Tile_i == 0 && Tile_j == 1 && BRAM_i == 1 && BRAM_j == 0) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
           
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
    if(Tile_i == 0 && Tile_j == 1 && BRAM_i == 1 && BRAM_j == 1) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
           
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end
	
	
	if(Tile_i == 1 && Tile_j == 0 && BRAM_i == 0 && BRAM_j == 0) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
           
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
    if(Tile_i == 1 && Tile_j == 0 && BRAM_i == 0 && BRAM_j == 1) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
            
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
    if(Tile_i == 1 && Tile_j == 0 && BRAM_i == 1 && BRAM_j == 0) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
           
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
    if(Tile_i == 1 && Tile_j == 0 && BRAM_i == 1 && BRAM_j == 1) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
           
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end
	
	
	if(Tile_i == 1 && Tile_j == 1 && BRAM_i == 0 && BRAM_j == 0) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
           
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
    if(Tile_i == 1 && Tile_j == 1 && BRAM_i == 0 && BRAM_j == 1) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
            
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
    if(Tile_i == 1 && Tile_j == 1 && BRAM_i == 1 && BRAM_j == 0) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
           
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end 
    if(Tile_i == 1 && Tile_j == 1 && BRAM_i == 1 && BRAM_j == 1) begin
        if(!reset) begin
            WEA = 1;
            for(k=15; k>=0; k=k-1) begin  
                DINA[k] = ram[k][ram_ptr];
            end
           
            ADDRA = ADDRA + 1;
            ram_ptr = ram_ptr + 1;
        end 
        else DINA = 0;
    end
	
end
initial
 
begin
//LENGTH = 16;
Tanh_In = 0;
Activation_Function = 0;
// 1001001010100100010010011011011
//    100101010010001001001101101111

// WEST_I = 'h33333333deadbeef00000000ffffffff00000003000000070000000b0000000f;
// WEST_I = 'h000000000000000000000000000000005555555555555555555555552548936f;
// instruction = 32'b000010_00001_00011_0000_0000_0000_0001;
reset = 0; 
start = 0;//0
mode = 0;
external = 1;

ram[0]  = 'h000010b3_00000001_00000000_00000000_00000000;
ram[1]  = 'h0000066f_00000002_00000000_00000000_00000000;
ram[2]  = 'h00000cec_000018b5_00000000_00000000_00000000;
ram[3]  = 'h000004D7_00007BE8_00000000_00010000_00000000;
ram[4]  = 'h000053F3_000044A7_00000000_00000000_00000000;
ram[5]  = 'hffffef4f_00000300_00000000_00000000_00000000;
ram[6] 	= 'h00123400_00ba2500_00000000_00000000_00000000;
ram[7] 	= 'h00965300_00003637_00000000_00020000_00000000;
ram[8] 	= 'hff753200_00123400_00000000_00000000_00000000;
ram[9] 	= 'h00325800_00965300_00000000_00000000_00000000;
ram[10]	= 'h00a25d00_00753200_00000000_00000000_00000000;
ram[11]	= 'h00d2b300_0000989A_00000000_00000000_00000000;
ram[12]	= 'hff501d00_ff354200_00000000_00000000_00000000;
ram[13]	= 'h00521000_00325700_00000000_00000000_00000000;
ram[14]	= 'h00862500_ffa25400_00000000_00000000_00000000;
ram[15]	= 'hffffff00_0000ABD5_00000000_00000000_00000000;
BRAM_i = 8'b0;
BRAM_j = 8'b0;
Tile_i = 8'b0;
Tile_j = 8'b0;
ADDRA = -1;
ram_ptr = 0;
#1610
ram[0]  = 'h00f41500_00ffff00_00000000_00000000_00000000;
ram[1]  = 'h00000000_00000021_00000000_00000000_00000000;
ram[2]  = 'h00456000_00003400_00000000_00000000_00000000;
ram[3]  = 'h00f41500_00ffff00_00000000_00000001_00000000;
ram[4]  = 'h00000000_00000560_00000000_00000000_00000000;
ram[5]  = 'h00000123_00201103_00000000_00000000_00000000;
ram[6] 	= 'h00325800_00000890_00000000_00000000_00000000;
ram[7] 	= 'h00000000_00ab0000_00000000_00000002_00000000;
ram[8] 	= 'h00000000_00521000_00000000_00000000_00000000;
ram[9] 	= 'h00000000_00000120_00000000_00000000_00000000;
ram[10]	= 'h00521000_00325700_00000000_00000000_00000000;
ram[11]	= 'h00000000_00000340_00000000_00000003_00000000;
ram[12]	= 'h00000000_00110000_00000000_00000000_00000000;
ram[13]	= 'h00000000_00000020_00000000_00000000_00000000;
ram[14]	= 'h00000000_00f6a000_00000000_00000000_00000000;
ram[15]	= 'h00000000_00001000_00000000_00000004_00000000;
BRAM_i = 8'b0;
BRAM_j = 8'b1;
Tile_i = 8'b0;
Tile_j = 8'b0;
ADDRA = -1;
ram_ptr = 0;
#1610
ram[0]  = 'h00000000_00000001_00000000_00000000_00000000;
ram[1]  = 'h00965300_00f41500_00000000_00020000_00000000;
ram[2]  = 'h00000000_00000002_00000000_00000000_00000000;
ram[3]  = 'h00000000_00654300_00000000_00000000_00000000;
ram[4]  = 'h00000000_00000003_00000000_00000000_00000000;
ram[5]  = 'hff501d00_ff354200_00000000_00000000_00000000;
ram[6] 	= 'h00000000_00000004_00000000_00000000_00000000;
ram[7] 	= 'h00000000_00000005_00000000_00000000_00000000;
ram[8] 	= 'h00f41500_00000006_00000000_00000000_00000000;
ram[9] 	= 'h00000000_00000007_00000000_00000000_00000000;
ram[10]	= 'h00000000_00000123_00000000_00000000_00000000;
ram[11]	= 'h00000000_00000008_00000000_00000000_00000000;
ram[12]	= 'h00000000_04560000_00000000_00000000_00000000;
ram[13]	= 'h00000000_00000009_00000000_00000000_00000000;
ram[14]	= 'h00000000_000abc00_00000000_00000000_00000000;
ram[15]	= 'h00000000_0000000a_00000000_00000000_00000000;
BRAM_i = 8'b1;
BRAM_j = 8'b0;
Tile_i = 8'b0;
Tile_j = 8'b0;
ADDRA = -1;
ram_ptr = 0;
#1610
ram[0]  = 'h00a25d00_00753200_00000000_00000000_00000000;
ram[1]  = 'h00000000_0000000b_00000000_00000000_00000000;
ram[2]  = 'h00123400_00ba2500_00000000_00000000_00000000;
ram[3]  = 'h000a2540_0000000c_00000000_00000005_00000000;
ram[4]  = 'h00000000_00000030_00000000_00000000_00000000;
ram[5]  = 'h00000000_0020000d_00000000_00000000_00000000;
ram[6] 	= 'h00000000_0000000e_00000000_00000000_00000000;
ram[7] 	= 'h00000000_0000000f_00000000_00000006_00000000;
ram[8] 	= 'h00000000_0000000a_00000000_00000000_00000000;
ram[9] 	= 'h00ba2500_ff862500_00000000_00000000_00000000;
ram[10]	= 'h00000000_00000001_00000000_00000000_00000000;
ram[11]	= 'h00000000_000008a0_00000000_00000007_00000000;
ram[12]	= 'h00000000_00000002_00000000_00000000_00000000;
ram[13]	= 'h00000000_00000440_00000000_00000000_00000000;
ram[14]	= 'h00000000_00000003_00000000_00000000_00000000;
ram[15]	= 'h00000000_00000550_00000000_00000008_00000000;
BRAM_i = 8'b1;
BRAM_j = 8'b1;
Tile_i = 8'b0;
Tile_j = 8'b0;
ADDRA = -1;
ram_ptr = 0;
#1610

ram[0]  = 'h00005678_12345678_00000000_00000000_00000000;
ram[1]  = 'h00354200_00d2b300_00000000_00000000_00000000;
ram[2]  = 'hff325700_00501d00_00000000_00000000_00000000;
ram[3]  = 'h00a25400_00654300_00000000_00010000_00000000;
ram[4]  = 'h00ba2500_ff862500_00000000_00000000_00000000;
ram[5]  = 'h00f41500_00ffff00_00000000_00000000_00000000;
ram[6] 	= 'h00123400_00ba2500_00000000_00000000_00000000;
ram[7] 	= 'h00965300_00f41500_00000000_00020000_00000000;
ram[8] 	= 'hff753200_00123400_00000000_00000000_00000000;
ram[9] 	= 'h00325800_00965300_00000000_00000000_00000000;
ram[10]	= 'h00a25d00_00753200_00000000_00000000_00000000;
ram[11]	= 'h00d2b300_00325800_00000000_00000000_00000000;
ram[12]	= 'hff501d00_ff354200_00000000_00000000_00000000;
ram[13]	= 'h00521000_00325700_00000000_00000000_00000000;
ram[14]	= 'h00862500_ffa25400_00000000_00000000_00000000;
ram[15]	= 'hffffff00_00521000_00000000_00000000_00000000;
BRAM_i = 8'b0;
BRAM_j = 8'b0;
Tile_i = 8'b0;
Tile_j = 8'b1;
ADDRA = -1;
ram_ptr = 0;
#1610
ram[0]  = 'h00f41500_00fabf00_00000000_00000000_00000000;
ram[1]  = 'h00000000_00000044_00000000_00000000_00000000;
ram[2]  = 'h00000000_00000050_00000000_00000000_00000000;
ram[3]  = 'h00f41500_00ffff00_00000000_00000000_00000000;
ram[4]  = 'h00000000_00000060_00000000_00000000_00000000;
ram[5]  = 'h00000000_00034000_00000000_00000000_00000000;
ram[6] 	= 'h00325800_00000070_00000000_00000000_00000000;
ram[7] 	= 'h00000000_00000080_00000000_00000002_00000000;
ram[8] 	= 'h00000000_00521000_00000000_00000000_00000000;
ram[9] 	= 'h00000000_00000090_00000000_00000000_00000000;
ram[10]	= 'h00521000_00325700_00000000_00000000_00000000;
ram[11]	= 'h00000000_00009800_00000000_00000003_00000000;
ram[12]	= 'h00000000_00000500_00000000_00000000_00000000;
ram[13]	= 'h00000000_000000a0_00000000_00000000_00000000;
ram[14]	= 'h00000000_000ab300_00000000_00000000_00000000;
ram[15]	= 'h00000000_00030020_00000000_00000004_00000000;
BRAM_i = 8'b0;
BRAM_j = 8'b1;
Tile_i = 8'b0;
Tile_j = 8'b1;
ADDRA = -1;
ram_ptr = 0;
#1610
ram[0]  = 'h00000000_00380000_00000000_00000000_00000000;
ram[1]  = 'h00965300_00f41500_00000000_00020000_00000000;
ram[2]  = 'h00000000_00000b00_00000000_00000000_00000000;
ram[3]  = 'h00000000_00654300_00000000_00000000_00000000;
ram[4]  = 'h00000000_00000c00_00000000_00000000_00000000;
ram[5]  = 'hff501d00_ff354200_00000000_00000000_00000000;
ram[6] 	= 'h00000000_00000d00_00000000_00000000_00000000;
ram[7] 	= 'h00000000_00000e00_00000000_00000000_00000000;
ram[8] 	= 'h00f41500_00000f00_00000000_00000000_00000000;
ram[9] 	= 'h00000000_00000a00_00000000_00000000_00000000;
ram[10]	= 'h00000000_00000100_00000000_00000000_00000000;
ram[11]	= 'h00000000_00098000_00000000_00000000_00000000;
ram[12]	= 'h00000000_00005500_00000000_00000000_00000000;
ram[13]	= 'h00000000_00030000_00000000_00000000_00000000;
ram[14]	= 'h00000000_00002010_00000000_00000000_00000000;
ram[15]	= 'h00000000_00504020_00000000_00000000_00000000;
BRAM_i = 8'b1;
BRAM_j = 8'b0;
Tile_i = 8'b0;
Tile_j = 8'b1;
ADDRA = -1;
ram_ptr = 0;
#1610
ram[0]  = 'h00a25d00_00753200_00000000_00000000_00000000;
ram[1]  = 'h00000000_00000200_00000000_00000000_00000000;
ram[2]  = 'h00123400_00ba2500_00000000_00000000_00000000;
ram[3]  = 'h000a2540_00000300_00000000_00000005_00000000;
ram[4]  = 'h00000000_00030000_00000000_00000000_00000000;
ram[5]  = 'h00000000_00000400_00000000_00000000_00000000;
ram[6] 	= 'h00000000_00000600_00000000_00000000_00000000;
ram[7] 	= 'h00000000_00000500_00000000_00000006_00000000;
ram[8] 	= 'h00000000_00007000_00000000_00000000_00000000;
ram[9] 	= 'h00ba2500_ff862500_00000000_00000000_00000000;
ram[10]	= 'h00000000_00008000_00000000_00000000_00000000;
ram[11]	= 'h00000000_00004040_00000000_00000007_00000000;
ram[12]	= 'h00000000_00000d30_00000000_00000000_00000000;
ram[13]	= 'h00000000_00ab0000_00000000_00000000_00000000;
ram[14]	= 'h00000000_00000200_00000000_00000000_00000000;
ram[15]	= 'h00000000_00098000_00000000_00000008_00000000;
BRAM_i = 8'b1;
BRAM_j = 8'b1;
Tile_i = 8'b0;
Tile_j = 8'b1;
ADDRA = -1;
ram_ptr = 0;
#1610


ram[0]  = 'h00005678_12345678_00000000_00000000_00000000;
ram[1]  = 'h00354200_00d2b300_00000000_00000000_00000000;
ram[2]  = 'hff325700_00501d00_00000000_00000000_00000000;
ram[3]  = 'h00a25400_00654300_00000000_00010000_00000000;
ram[4]  = 'h00ba2500_ff862500_00000000_00000000_00000000;
ram[5]  = 'h00f41500_00ffff00_00000000_00000000_00000000;
ram[6] 	= 'h00123400_00ba2500_00000000_00000000_00000000;
ram[7] 	= 'h00965300_00f41500_00000000_00020000_00000000;
ram[8] 	= 'hff753200_00123400_00000000_00000000_00000000;
ram[9] 	= 'h00325800_00965300_00000000_00000000_00000000;
ram[10]	= 'h00a25d00_00753200_00000000_00000000_00000000;
ram[11]	= 'h00d2b300_00325800_00000000_00000000_00000000;
ram[12]	= 'hff501d00_ff354200_00000000_00000000_00000000;
ram[13]	= 'h00521000_00325700_00000000_00000000_00000000;
ram[14]	= 'h00862500_ffa25400_00000000_00000000_00000000;
ram[15]	= 'hffffff00_00521000_00000000_00000000_00000000;
BRAM_i = 8'b0;
BRAM_j = 8'b0;
Tile_i = 8'b1;
Tile_j = 8'b0;
ADDRA = -1;
ram_ptr = 0;
#1610
ram[0]  = 'h00f41500_00ffff00_00000000_00000000_00000000;
ram[1]  = 'h00000000_00009000_00000000_00000000_00000000;
ram[2]  = 'h00000000_0000a000_00000000_00000000_00000000;
ram[3]  = 'h00f41500_00ffff00_00000000_00000000_00000000;
ram[4]  = 'h00000000_0000b000_00000000_00000000_00000000;
ram[5]  = 'h00000000_0000c000_00000000_00000000_00000000;
ram[6] 	= 'h00325800_00520000_00000000_00000000_00000000;
ram[7] 	= 'h00000000_00000050_00000000_00000002_00000000;
ram[8] 	= 'h00000000_00521000_00000000_00000000_00000000;
ram[9] 	= 'h00000000_0000d000_00000000_00000000_00000000;
ram[10]	= 'h00521000_00325700_00000000_00000000_00000000;
ram[11]	= 'h00000000_0000e000_00000000_00000003_00000000;
ram[12]	= 'h00000000_00066000_00000000_00000000_00000000;
ram[13]	= 'h00000000_00000050_00000000_00000000_00000000;
ram[14]	= 'h00000000_00043000_00000000_00000000_00000000;
ram[15]	= 'h00000000_00000770_00000000_00000004_00000000;
BRAM_i = 8'b0;
BRAM_j = 8'b1;
Tile_i = 8'b1;
Tile_j = 8'b0;
ADDRA = -1;
ram_ptr = 0;
#1610
ram[0]  = 'h00000000_000f0000_00000000_00000000_00000000;
ram[1]  = 'h00965300_00f41500_00000000_00020000_00000000;
ram[2]  = 'h00000000_000a0000_00000000_00000000_00000000;
ram[3]  = 'h00000000_00654300_00000000_00000000_00000000;
ram[4]  = 'h00000000_00010000_00000000_00000000_00000000;
ram[5]  = 'hff501d00_ff354200_00000000_00000000_00000000;
ram[6] 	= 'h00000000_00020000_00000000_00000000_00000000;
ram[7] 	= 'h00000000_00030000_00000000_00000000_00000000;
ram[8] 	= 'h00f41500_00040000_00000000_00000000_00000000;
ram[9] 	= 'h00000000_00050000_00000000_00000000_00000000;
ram[10]	= 'h00000000_00230000_00000000_00000000_00000000;
ram[11]	= 'h00000000_00060000_00000000_00000000_00000000;
ram[12]	= 'h00000000_00000608_00000000_00000000_00000000;
ram[13]	= 'h00000000_00200400_00000000_00000000_00000000;
ram[14]	= 'h00000000_0a0b00c0_00000000_00000000_00000000;
ram[15]	= 'h00000000_0000a050_00000000_00000000_00000000;
BRAM_i = 8'b1;
BRAM_j = 8'b0;
Tile_i = 8'b1;
Tile_j = 8'b0;
ADDRA = -1;
ram_ptr = 0;
#1610
ram[0]  = 'h00a25d00_00753200_00000000_00000000_00000000;
ram[1]  = 'h00000000_00007000_00000000_00000000_00000000;
ram[2]  = 'h00123400_00ba2500_00000000_00000000_00000000;
ram[3]  = 'h000a2540_00080000_00000000_00000005_00000000;
ram[4]  = 'h00000000_00b00000_00000000_00000000_00000000;
ram[5]  = 'h00000000_00090000_00000000_00000000_00000000;
ram[6] 	= 'h00000000_000000a0_00000000_00000000_00000000;
ram[7] 	= 'h00000000_000b0000_00000000_00000006_00000000;
ram[8] 	= 'h00000000_000c0000_00000000_00000000_00000000;
ram[9] 	= 'h00ba2500_ff862500_00000000_00000000_00000000;
ram[10]	= 'h00000000_000d0000_00000000_00000000_00000000;
ram[11]	= 'h00000000_0c000000_00000000_00000007_00000000;
ram[12]	= 'h00000000_00000c00_00000000_00000000_00000000;
ram[13]	= 'h00000000_0200b000_00000000_00000000_00000000;
ram[14]	= 'h00000000_00d00600_00000000_00000000_00000000;
ram[15]	= 'h00000000_00da0400_00000000_00000008_00000000;
BRAM_i = 8'b1;
BRAM_j = 8'b1;
Tile_i = 8'b1;
Tile_j = 8'b0;
ADDRA = -1;
ram_ptr = 0;
#1610

ram[0]  = 'h00005678_12345678_00000000_00000000_00000000;
ram[1]  = 'h00354200_00d2b300_00000000_00000000_00000000;
ram[2]  = 'hff325700_00501d00_00000000_00000000_00000000;
ram[3]  = 'h00a25400_00654300_00000000_00010000_00000000;
ram[4]  = 'h00ba2500_ff862500_00000000_00000000_00000000;
ram[5]  = 'h00f41500_00ffff00_00000000_00000000_00000000;
ram[6] 	= 'h00123400_00ba2500_00000000_00000000_00000000;
ram[7] 	= 'h00965300_00f41500_00000000_00020000_00000000;
ram[8] 	= 'hff753200_00123400_00000000_00000000_00000000;
ram[9] 	= 'h00325800_00945400_00000000_00000000_00000000;
ram[10]	= 'h00a25d00_00743200_00000000_00000000_00000000;
ram[11]	= 'h00d2b300_00323400_00000000_00000000_00000000;
ram[12]	= 'hff501d00_ff354200_00000000_00000000_00000000;
ram[13]	= 'h00521000_00323700_00000000_00000000_00000000;
ram[14]	= 'h00862500_ffa25400_00000000_00000000_00000000;
ram[15]	= 'hffffff00_00523000_00000000_00000000_00000000;
BRAM_i = 8'b0;
BRAM_j = 8'b0;
Tile_i = 8'b1;
Tile_j = 8'b1;
ADDRA = -1;
ram_ptr = 0;
#1610
ram[0]  = 'h00f41500_00ffff00_00000000_00000000_00000000;
ram[1]  = 'h00000000_000e0000_00000000_00000000_00000000;
ram[2]  = 'h00000000_00000ff0_00000000_00000000_00000000;
ram[3]  = 'h00f41500_00fffd00_00000000_00000000_00000000;
ram[4]  = 'h00000000_000a0000_00000000_00000000_00000000;
ram[5]  = 'h00000000_0000d000_00000000_00000000_00000000;
ram[6] 	= 'h00325800_00a00000_00000000_00000000_00000000;
ram[7] 	= 'h00000000_00100000_00000000_00000002_00000000;
ram[8] 	= 'h00000000_00521000_00000000_00000000_00000000;
ram[9] 	= 'h00000000_00200000_00000000_00000000_00000000;
ram[10]	= 'h00521000_00325700_00000000_00000000_00000000;
ram[11]	= 'h00000000_00300000_00000000_00000003_00000000;
ram[12]	= 'h00000000_00b000c0_00000000_00000000_00000000;
ram[13]	= 'h00000000_00000a00_00000000_00000000_00000000;
ram[14]	= 'h00000000_00b00000_00000000_00000000_00000000;
ram[15]	= 'h00000000_000d0c00_00000000_00000004_00000000;
BRAM_i = 8'b0;
BRAM_j = 8'b1;
Tile_i = 8'b1;
Tile_j = 8'b1;
ADDRA = -1;
ram_ptr = 0;
#1610
ram[0]  = 'h00000000_00300000_00000000_00000000_00000000;
ram[1]  = 'h00965300_00f41500_00000000_00020000_00000000;
ram[2]  = 'h00000000_00040000_00000000_00000000_00000000;
ram[3]  = 'h00000000_00654300_00000000_00000000_00000000;
ram[4]  = 'h00000000_00000000_00000000_00000000_00000000;
ram[5]  = 'hff501d00_ff354200_00000000_00000000_00000000;
ram[6] 	= 'h00000000_00500000_00000000_00000000_00000000;
ram[7] 	= 'h00000000_00600000_00000000_00000000_00000000;
ram[8] 	= 'h00f41500_00010000_00000000_00000000_00000000;
ram[9] 	= 'h00000000_00600000_00000000_00000000_00000000;
ram[10]	= 'h00000000_00070000_00000000_00000000_00000000;
ram[11]	= 'h00000000_00010200_00000000_00000000_00000000;
ram[12]	= 'h00000000_00000003_00000000_00000000_00000000;
ram[13]	= 'h00000000_00305000_00000000_00000000_00000000;
ram[14]	= 'h00000000_00200060_00000000_00000000_00000000;
ram[15]	= 'h00000000_00045400_00000000_00000000_00000000;
BRAM_i = 8'b1;
BRAM_j = 8'b0;
Tile_i = 8'b1;
Tile_j = 8'b1;
ADDRA = -1;
ram_ptr = 0;
#1610
ram[0]  = 'h00a25d00_00753200_00000000_00000000_00000000;
ram[1]  = 'h00000000_00800000_00000000_00000000_00000000;
ram[2]  = 'h00123400_00ba2500_00000000_00000000_00000000;
ram[3]  = 'h000a2540_00090000_00000000_00000005_00000000;
ram[4]  = 'h00000000_00a00000_00000000_00000000_00000000;
ram[5]  = 'h00000000_00b00000_00000000_00000000_00000000;
ram[6] 	= 'h00000000_00007000_00000000_00000000_00000000;
ram[7] 	= 'h00000000_00c00000_00000000_00000006_00000000;
ram[8] 	= 'h00000000_00d00000_00000000_00000000_00000000;
ram[9] 	= 'h00ba2500_ff862700_00000000_00000000_00000000;
ram[10]	= 'h00000000_00c000d0_00000000_00000000_00000000;
ram[11]	= 'h00000000_0000c000_00000000_00000007_00000000;
ram[12]	= 'h00000000_0d0900e0_00000000_00000000_00000000;
ram[13]	= 'h00000000_00b00a00_00000000_00000000_00000000;
ram[14]	= 'h00000000_00080080_00000000_00000000_00000000;
ram[15]	= 'h00000000_00a0b090_00000000_00000008_00000000;
BRAM_i = 8'b1;
BRAM_j = 8'b1;
Tile_i = 8'b1;
Tile_j = 8'b1;
ADDRA = -1;
ram_ptr = 0;
#1610


DINA = 0;
#10
external = 0;
#10000
reset = 1;//1 
#2000

// // DIN = 16'hFFFF;
// instruction = (2<<26) + (1<<21) + (3<<16) + (4<<11);
// start = 1;
// #124
// start = 0;//1
#1000

Activation_Function = 2'b00;
Tanh_In = 0;
//////////////////////////////////////////////////////
//instruction = (5<<26) + (1<<21) + (3<<16) + (1<<11);
//instruction = (0<<26) + (1<<21) + (3<<16) + (4<<11);
//start = 1;
//#100 start = 0;
//#1000
instruction = (5<<26) + (1<<21) + (3<<16) + (2<<11);
start = 1;
#100 start = 0;
//#1000
//instruction = (7<<26) + (3<<21) + (3<<16) + (1<<11);
//start = 1;
//#100 start = 0;
//////////////////////////////////////////////////
// #10000
// //////////////////////////////////////////////////////
// instruction = (2<<26) + (2<<21) + (3<<16) + (4<<11);
// start = 1;
// #100 start = 0;
// ////////////////////////////////////////////////////
// ////////////////////////////////////////////////////
//#10000
//Activation_Function = 2;
//Tanh_In = 1;
// //////////////////////////////////////////////////////
// //////////////////////////////////////////////////////
// instruction = (8<<26) + (1<<21) + (1<<16) + (0<<11);
// start = 1;
// #10 start = 0;//1
// //////////////////////////////////////////////////////
// #10000
// //////////////////////////////////////////////////////
// instruction = (7<<26) + (1<<21) + (1<<16) + (0<<11);
// start = 1;
// #10 start = 0;//1
// // //////////////////////////////////////////////////////






// #1000
// instruction = (7<<26) + (0<<21) + (0<<16) + (0<<11);
// #100
// start = 1;
// #124
// start = 0;//1
// #1000
// start = 1;
// #124
// start = 0;//1

// reset = 0;
// #1000
// reset = 1;
// #1000
// start = 1;
// #113
// start = 0;//1
// // mode = 1;
// // #100
// start = 1;
// #10
// start = 0;
// // DIN = 16'hFFFF;
// instruction = 32'h14221800;
// start = 1;
// #10 
// start = 0;//1
// #1000
// start = 1;
// #10 
// start = 0;//1
// #1000
// start = 1;
// #10 
// start = 0;//1

// instruction = 32'b000100_00001_00011_0000_0000_0000_0000;
// #30000
// start = 1;
// #10
// start = 0;
// #200000
// LENGTH = 16;
// reset = 0;
// start = 0;
// block_addr = 0;
// reg_addr = 0;
// #30000 
// reg_addr = 'h10;
// block_addr = 0;
// reset = 1;
// start = 1;
// #20000
// start = 0;


end

endmodule